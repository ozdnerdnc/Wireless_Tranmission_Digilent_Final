----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 26.04.2018 19:34:07
-- Design Name: 
-- Module Name: ROM - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ROM is
    Port ( a : in STD_LOGIC_VECTOR (13 downto 0);
           spo : out STD_LOGIC_VECTOR ( 2 downto 0)
           );
end ROM;

architecture Behavioral of ROM is
-- Block ROM 
type vector_array is ARRAY (0 to 10799) of std_logic_vector (2 downto 0); 
-- Initialization code taken from .coe file
signal memory: vector_array := ("111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"000",
"000",
"111",
"111",
"000",
"000",
"111",
"000",
"000",
"111",
"111",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"000",
"110",
"000",
"111",
"111",
"000",
"110",
"000",
"111",
"000",
"110",
"110",
"000",
"001",
"111",
"111",
"001",
"110",
"111",
"000",
"000",
"111",
"000",
"111",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"000",
"111",
"000",
"110",
"110",
"000",
"001",
"110",
"110",
"110",
"000",
"110",
"110",
"110",
"000",
"110",
"110",
"111",
"000",
"110",
"111",
"000",
"000",
"111",
"001",
"001",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"000",
"110",
"110",
"110",
"110",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"110",
"110",
"110",
"111",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"000",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"001",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"001",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"001",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"110",
"110",
"110",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"001",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"001",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"001",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"001",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"110",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"000",
"000",
"000",
"110",
"110",
"110",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"110",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"001",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"001",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"111",
"001",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"001",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"000",
"100",
"100",
"100",
"000",
"000",
"111",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"100",
"100",
"100",
"100",
"000",
"000",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"100",
"100",
"100",
"100",
"100",
"000",
"000",
"100",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"000",
"100",
"100",
"100",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"100",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"001",
"000",
"110",
"110",
"110",
"110",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"000",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"000",
"000",
"100",
"111",
"111",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"001",
"000",
"000",
"110",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"000",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"011",
"000",
"100",
"100",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"000",
"000",
"100",
"100",
"100",
"100",
"100",
"000",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"000",
"100",
"100",
"100",
"100",
"000",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"000",
"110",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"100",
"100",
"100",
"100",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"000",
"110",
"110",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"000",
"000",
"100",
"100",
"000",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"000",
"000",
"100",
"100",
"100",
"100",
"000",
"110",
"110",
"110",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"100",
"000",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"011",
"000",
"100",
"100",
"100",
"100",
"000",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"110",
"110",
"110",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"000",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"111",
"000",
"100",
"100",
"100",
"100",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"000",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"000",
"111",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"000",
"100",
"100",
"100",
"100",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"010",
"010",
"010",
"010",
"010",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"000",
"000",
"100",
"100",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"010",
"000",
"010",
"000",
"110",
"110",
"110",
"000",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"111",
"111",
"000",
"100",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"010",
"000",
"010",
"000",
"110",
"110",
"110",
"000",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"111",
"111",
"000",
"111",
"111",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"010",
"010",
"010",
"010",
"010",
"000",
"110",
"110",
"000",
"000",
"110",
"110",
"000",
"111",
"000",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"010",
"000",
"010",
"010",
"000",
"110",
"000",
"000",
"000",
"110",
"110",
"000",
"110",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"111",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"101",
"010",
"010",
"010",
"000",
"010",
"010",
"000",
"010",
"010",
"111",
"001",
"110",
"000",
"111",
"111",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"101",
"010",
"010",
"010",
"110",
"010",
"010",
"000",
"010",
"000",
"000",
"111",
"000",
"111",
"111",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"010",
"010",
"010",
"111",
"010",
"010",
"010",
"010",
"000",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"010",
"010",
"010",
"110",
"010",
"010",
"111",
"010",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"111",
"000",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"010",
"010",
"010",
"110",
"010",
"010",
"111",
"010",
"000",
"111",
"111",
"111",
"111",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"111",
"000",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"000",
"000",
"000",
"010",
"010",
"010",
"110",
"010",
"010",
"110",
"010",
"000",
"111",
"111",
"111",
"111",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"000",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"111",
"111",
"000",
"000",
"000",
"000",
"010",
"010",
"010",
"110",
"010",
"010",
"110",
"010",
"000",
"111",
"111",
"111",
"111",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"001",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"010",
"010",
"010",
"110",
"010",
"010",
"110",
"010",
"000",
"111",
"111",
"111",
"111",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"111",
"110",
"110",
"001",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"010",
"010",
"010",
"110",
"010",
"010",
"110",
"010",
"000",
"111",
"111",
"111",
"111",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"111",
"111",
"110",
"111",
"000",
"001",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"010",
"010",
"010",
"110",
"010",
"010",
"010",
"010",
"010",
"111",
"111",
"111",
"111",
"111",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"000",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"010",
"010",
"010",
"110",
"010",
"010",
"000",
"010",
"010",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"000",
"000",
"000",
"110",
"000",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"010",
"010",
"010",
"110",
"010",
"010",
"000",
"010",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"000",
"000",
"000",
"000",
"000",
"110",
"110",
"000",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"010",
"010",
"010",
"110",
"010",
"010",
"010",
"010",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"100",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"110",
"110",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"010",
"010",
"010",
"110",
"010",
"010",
"110",
"010",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"000",
"001",
"001",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"010",
"010",
"010",
"110",
"010",
"010",
"110",
"010",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"010",
"010",
"010",
"111",
"010",
"010",
"111",
"010",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"010",
"010",
"010",
"110",
"010",
"010",
"110",
"010",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"110",
"010",
"010",
"010",
"010",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"110",
"010",
"010",
"110",
"010",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"010",
"010",
"110",
"010",
"010",
"110",
"010",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"111",
"010",
"010",
"110",
"010",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"110",
"010",
"010",
"010",
"110",
"111",
"101",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"110",
"110",
"010",
"010",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"010",
"110",
"010",
"010",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"110",
"010",
"010",
"010",
"110",
"010",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"000",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"110",
"110",
"010",
"010",
"110",
"010",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"001",
"000",
"110",
"110",
"001",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"010",
"010",
"010",
"110",
"010",
"010",
"110",
"010",
"111",
"101",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"001",
"001",
"000",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"010",
"010",
"010",
"110",
"010",
"010",
"110",
"010",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"110",
"000",
"111",
"111",
"000",
"000",
"111",
"111",
"000",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"010",
"010",
"010",
"110",
"010",
"010",
"111",
"010",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"001",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"000",
"111",
"111",
"000",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"111",
"000",
"000",
"000",
"000",
"010",
"010",
"010",
"111",
"010",
"010",
"110",
"010",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"000",
"111",
"111",
"000",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"111",
"111",
"111",
"000",
"000",
"000",
"010",
"010",
"010",
"111",
"010",
"010",
"111",
"110",
"111",
"101",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"010",
"010",
"111",
"010",
"010",
"110",
"010",
"111",
"101",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"001",
"000",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"110",
"000",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"010",
"010",
"111",
"010",
"010",
"010",
"110",
"010",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"010",
"010",
"110",
"110",
"010",
"010",
"010",
"010",
"010",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"000",
"010",
"010",
"110",
"111",
"010",
"010",
"010",
"010",
"111",
"101",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"010",
"111",
"010",
"010",
"010",
"010",
"010",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"111",
"010",
"010",
"010",
"010",
"010",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"010",
"010",
"111",
"010",
"010",
"010",
"010",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"110",
"110",
"010",
"010",
"010",
"110",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"111",
"010",
"010",
"010",
"010",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"010",
"010",
"110",
"111",
"010",
"010",
"010",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"010",
"010",
"110",
"110",
"010",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"000",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"000",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111",
"111"




 );


begin
      
spo<=memory(conv_integer(a)) ; 	

	 

end Behavioral;
